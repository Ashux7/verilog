module test;
initial begin
$display("Heloo");
$finish;
end
endmodule

