`timescale 1ps/1ps

module q2;

    reg A

endmodule