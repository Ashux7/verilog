`timescale 1ps/1ps
module OR (
    input A,
    input B,
    output Y
);
    assign Y = A|B;
endmodule
